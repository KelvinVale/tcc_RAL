O que tem para fazer :


	agents:
		-agent_in
			.interfacee			pendente
			.transaction		pendente
			.sequence			pendente
			.sequencer			pendente
			.driver				pendente
			.monitor			pendente
			.montar_agent		pendente

		-agent_out
			.interfacee			pendente
			.transaction		pendente
			.driver				pendente
			.monitor			pendente
			.montar_agent		pendente

	scoreboard:
		-refmods
			.refmod.c				pendente
			.refmod.sv				pendente
		-comparador					pendente
		-montar_scoreboard			pendente

	env:
		-agents						pendente
		-scoreboard					pendente
		-cobertura					pendente
		-montar_env					pendente

	teste:
		-env 						pendente
		-montar_teste				pendente //Ativar a sequência !!!!

	top:
		-dut						pendente
		-montar_top					pendente




	Mudar arquivo 'pkg' 			pendente

	Mudar Makefile 					pendente


